--FOR EP3C16Q240C8
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use ieee.numeric_std.all;

entity OLED128x32 is
port(    	      	                                      --���}����   
        ck, nReset  :in std_logic;                     --�_����J(149) & RESET���s(145) 
        TSL2561_sda : INOUT  STD_LOGIC;                 --TSL2561 IIC SDA()
        TSL2561_scl : INOUT  STD_LOGIC;                 --TSL2561 IIC SCL()                  

		RSin : in std_logic;				--RS232
		RSout : out std_logic;
		
        SD178_sda  : INOUT  STD_LOGIC;                  --SD178B IIC SDA() 
        SD178_scl  : INOUT  STD_LOGIC;                  --SD178B IICSCL()     
        SD178_nrst : buffer    STD_LOGIC;                  --SD178B nRESET () 
        
        out_g		  :buffer std_logic_vector(7 downto 0);
		out_r			  :buffer std_logic_vector(7 downto 0);
		com		  :buffer std_logic_vector(7 downto 0); 
	
        SHT11_PIN : inout  STD_LOGIC;                   -- DHT11 PIN 

        sw    : IN std_logic_vector(7 downto 0);    --DIP SW()
        ki   : IN std_logic_vector(3 downto 0);        --BUTTON ()               
        ko  : buffer  std_logic_vector(3 downto 0);  
       -- debug  : OUT    STD_LOGIC;  
        	
        segout  :buffer std_logic_vector(7 downto 0);      --����C�q��ܾ���Ƹ}()
        segout_2:buffer std_logic_vector(7 downto 0);      --�k��C�q��ܾ���Ƹ}()       	        	        	
        seg_scan:buffer std_logic_vector(7 downto 0);          --�k��C�q��ܾ����y�}()           
                
        BL,RES,CS,DC,SDA,SCL : OUT    STD_LOGIC;        --LCD
        
        LED:buffer std_logic_vector(15 downto 0);
        LED_R,LED_G,LED_Y,buzzer:buffer std_logic;
        LED_RGB:buffer std_logic_vector(2 downto 0);
        
       -- PWM1,PWM2:out std_logic;
        
        motor_out1,motor_out2,motor_pwm1 : OUT    STD_LOGIC;
        motor_out3,motor_out4,motor_pwm2 : OUT    STD_LOGIC
         
    );
end OLED128x32;
architecture beh of OLED128x32 is

component i2c_master is
  GENERIC(
    input_clk : INTEGER := 50_000_000; --input clock speed from user logic in Hz
    bus_clk   : INTEGER := 100_000);   --speed the i2c bus (scl) will run at in Hz
  PORT(
    clk       : IN     STD_LOGIC;                    --system clock
    reset_n   : IN     STD_LOGIC;                    --active low reset
    ena       : IN     STD_LOGIC;                    --latch in command
    addr      : IN     STD_LOGIC_VECTOR(6 DOWNTO 0); --address of target slave
    rw        : IN     STD_LOGIC;                    --'0' is write, '1' is read
    data_wr   : IN     STD_LOGIC_VECTOR(7 DOWNTO 0); --data to write to slave
    busy      : OUT    STD_LOGIC;                    --indicates transaction in progress
    data_rd   : OUT    STD_LOGIC_VECTOR(7 DOWNTO 0); --data read from slave
    ack_error : BUFFER STD_LOGIC;                    --flag if improper acknowledge from slave
    sda       : INOUT  STD_LOGIC;                    --serial data output of i2c bus
    scl       : INOUT  STD_LOGIC);                   --serial clock output of i2c bus
end component i2c_master; 

component TSL2561 is 
port(
	  clk_50M:in std_logic;
     nrst:in std_logic;

     sda       : INOUT  STD_LOGIC;                   --TSL2561 IIC SDA(161)
     scl       : INOUT  STD_LOGIC;                   --TSL2561 IIC SCL(160)                                                             
     
     TSL2561_data : OUT  std_logic_vector(14 downto 0)

     );
end component TSL2561;

component DHT11 is 
port(
	   clk_50M:in std_logic;
     nrst:in std_logic;
     dat_bus: inout std_logic;
     HU, TE:out std_logic_vector(7 downto 0);        --????, ????
     error: out std_logic
     
     );
end component DHT11;

component cmd_rom is
   port(    
        address   : IN std_logic_vector(15 downto 0); 
        data_out  : OUT std_logic_vector(7 downto 0); 
        DC_data   : OUT std_logic   
       );
end component cmd_rom;

--component raminfr is
--generic ( 
--          bits : integer := 6;                -- number of bits per RAM word
--          addr_bits : integer := 15);         -- 2^addr_bits = number of words in RAM
--
--port (clk : in std_logic;
--       we : in std_logic;
--        a : in std_logic_vector(addr_bits-1 downto 0);
--       di : in std_logic_vector(bits-1 downto 0);
--       do : out std_logic_vector(bits-1 downto 0));
--end component raminfr;   
            
type State_type3 is (sd178_init, event_check, sd178_send , sd178_d1, sd178_d2, sd178_d3, sd178_d4, sd178_d5, sd178_delay1,sd178_delay2, sd178_set_ch,sd178_play1,sd178_play2);
SIGNAL  sd178State  : State_type3; 

type State_type4 is (event_check, s0, s1, s2, s3, s4, button1_process, button2_process, button3_process, button4_process, button5_process);
SIGNAL  Main_State  : State_type4;
--LCD NUMBER DATA
type oled_num_16x16 is array (48 to 122,0 to 15) of std_logic_vector(0 to 15);       --ASCII 0~z
constant num_table1:oled_num_16x16:=
(   
   (
   	X"0000",	X"0000",	X"03e0",	X"1c18",	X"300c",	X"300c",	X"7006",	X"6006",--0
   	X"6006",	X"6006",	X"300c",	X"300c",	X"1818",	X"07f0",	X"0000",	X"0000"
   ),
   (
	   X"0000",	X"0000",	X"0080",	X"0f80",	X"0180",	X"0180",	X"0180",	X"0180",--1
	   X"0180",	X"0180",	X"0180",	X"0180",	X"0180",	X"0ff0",	X"0000",	X"0000"  
   ),   
   (   
	  X"0000",	X"0000",	X"07c0",	X"1870",	X"2018",	X"4018",	X"0018",	X"0010",--2
	  X"0030",	X"00c0",	X"0100",	X"0600",	X"0806",	X"7ffc",	X"0000",	X"0000"   
   ),
   (
   	X"0000",	X"0000",	X"07e0",	X"1830",	X"2018",	X"0010",	X"0020",	X"01e0",--3
   	X"0638",	X"001c",	X"000c",	X"0008",	X"0010",	X"3fe0",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"0010",	X"0070",	X"00b0",	X"0130",	X"0230",	X"0c30",--4
   	X"1830",	X"2030",	X"7ffe",	X"0030",	X"0030",	X"0030",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"03fc",	X"0600",	X"0400",	X"0c00",	X"1fe0",	X"0070",--5
   	X"0018",	X"000c",	X"000c",	X"0008",	X"0010",	X"3fe0",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"003c",	X"03c0",	X"0600",	X"1800",	X"31c0",	X"3e38",--6
   	X"700c",	X"600c",	X"2006",	X"3004",	X"1808",	X"07f0",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"1ffc",	X"100c",	X"2008",	X"0018",	X"0010",	X"0030",--7
   	X"0060",	X"0060",	X"00c0",	X"0080",	X"0180",	X"0300",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"07e0",	X"1818",	X"3008",	X"3018",	X"1c30",	X"07c0",--8
   	X"06e0",	X"1838",	X"300c",	X"3006",	X"300c",	X"0ff0",	X"0000",	X"0000"
   ),
   (
   	X"0000",	X"0000",	X"07c0",	X"1830",	X"300c",	X"200c",	X"700c",	X"300c",--9
   	X"180c",	X"07fc",	X"0018",	X"0030",	X"00c0",	X"3f00",	X"0000",	X"0000"
   ),
   
(
	 
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"03c0",	x"0380",
	x"0000",	x"0000",	x"0000",	x"0000",	x"03c0",	x"0380",	x"0000",	x"0000"
),

(
	 
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"03c0",	x"0380",
	x"0000",	x"0000",	x"0000",	x"0100",	x"03c0",	x"00c0",	x"0080",	x"0300"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0000",	x"0006",	x"0038",	x"00c0",	x"0700",	x"1800",
	x"3000",	x"0e00",	x"0180",	x"0060",	x"001c",	x"0002",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"7ffe",	x"0000",
	x"0000",	x"7ffe",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0000",	x"3000",	x"0c00",	x"0300",	x"00e0",	x"0018",
	x"000c",	x"0070",	x"0180",	x"0600",	x"3800",	x"0000",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"1ff8",	x"200c",	x"700e",	x"380c",	x"0038",	x"00c0",
	x"0180",	x"0100",	x"0100",	x"0000",	x"0780",	x"0380",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0ff0",	x"180c",	x"3004",	x"63f2",	x"6632",	x"6662",
	x"6c64",	x"6c64",	x"6cc8",	x"6772",	x"3004",	x"1808",	x"07f0",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0180",	x"01c0",	x"02c0",	x"04c0",	x"04e0",	x"0460",
	x"0870",	x"0fb0",	x"1038",	x"1018",	x"2018",	x"787e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ff0",	x"181c",	x"180c",	x"181c",	x"1838",	x"1fe0",
	x"181c",	x"1806",	x"1806",	x"180e",	x"181c",	x"7fe0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0ffc",	x"1804",	x"3002",	x"7000",	x"6000",	x"6000",
	x"6000",	x"6000",	x"7002",	x"3804",	x"1c08",	x"03f0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3fc0",	x"1838",	x"180c",	x"180e",	x"1806",	x"1806",
	x"1806",	x"180e",	x"180c",	x"1818",	x"1860",	x"7f80",	x"0000",	x"0000"
),                                                                                            
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ffc",	x"180c",	x"1804",	x"1860",	x"1860",	x"1fe0",
	x"1860",	x"1860",	x"1802",	x"1806",	x"180c",	x"7ffc",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ffc",	x"180c",	x"1804",	x"1860",	x"1860",	x"1fe0",
	x"1860",	x"1860",	x"1800",	x"1800",	x"1800",	x"7e00",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0ffc",	x"180c",	x"3004",	x"7000",	x"6000",	x"6000",
	x"607e",	x"6018",	x"7018",	x"3018",	x"1818",	x"07e0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3c3c",	x"181c",	x"181c",	x"181c",	x"181c",	x"1ffc",
	x"181c",	x"181c",	x"181c",	x"181c",	x"181c",	x"7e7e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"07e0",	x"0180",	x"0180",	x"0180",	x"0180",	x"0180",
	x"0180",	x"0180",	x"0180",	x"0180",	x"0180",	x"0ff0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"03f8",	x"00e0",	x"00e0",	x"00e0",	x"00e0",	x"00e0",
	x"00e0",	x"00e0",	x"00e0",	x"00e0",	x"38c0",	x"1f00",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3c38",	x"3820",	x"3840",	x"3880",	x"3900",	x"3f00",
	x"3980",	x"38c0",	x"38e0",	x"3870",	x"3838",	x"7e7e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3e00",	x"1800",	x"1800",	x"1800",	x"1800",	x"1800",
	x"1800",	x"1800",	x"1800",	x"1802",	x"180e",	x"7ffc",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"783c",	x"383c",	x"383c",	x"2c5c",	x"2c5c",	x"2c5c",
	x"269c",	x"269c",	x"239c",	x"231c",	x"231c",	x"f83e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"380c",	x"1c08",	x"1608",	x"1708",	x"1388",	x"1188",
	x"10c8",	x"1068",	x"1038",	x"1038",	x"1018",	x"7c08",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0ff0",	x"1818",	x"300c",	x"700e",	x"6006",	x"6006",
	x"6006",	x"6006",	x"700c",	x"300c",	x"1810",	x"07e0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ff8",	x"180c",	x"1806",	x"1806",	x"180e",	x"1878",
	x"1f80",	x"1800",	x"1800",	x"1800",	x"1800",	x"7e00",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0ff0",	x"181c",	x"300c",	x"700e",	x"6006",	x"6006",
	x"6006",	x"6006",	x"770e",	x"38cc",	x"1878",	x"07e0",	x"003e",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ff0",	x"381c",	x"380e",	x"380e",	x"381c",	x"3fe0",
	x"39c0",	x"38e0",	x"3860",	x"3830",	x"3818",	x"7e1e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"1ffc",	x"300c",	x"3006",	x"3800",	x"1e00",	x"07e0",
	x"007c",	x"000e",	x"4006",	x"2006",	x"380c",	x"17f0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"7ffe",	x"6186",	x"4182",	x"0180",	x"0180",	x"0180",
	x"0180",	x"0180",	x"0180",	x"0180",	x"0180",	x"0ff0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3c0c",	x"180c",	x"180c",	x"180c",	x"180c",	x"180c",
	x"180c",	x"180c",	x"180c",	x"1808",	x"1c18",	x"07e0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3c1c",	x"1c08",	x"1c08",	x"0c10",	x"0e10",	x"0620",
	x"0720",	x"0740",	x"0340",	x"0380",	x"0180",	x"0100",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"71c6",	x"30c4",	x"30c4",	x"39cc",	x"19c8",	x"1968",
	x"1a68",	x"0e70",	x"0e70",	x"0c30",	x"0c20",	x"0420",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"1c1c",	x"0c10",	x"0e20",	x"0740",	x"0380",	x"0180",
	x"02c0",	x"02e0",	x"0460",	x"0830",	x"1038",	x"787e",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"380c",	x"1808",	x"1c10",	x"0e30",	x"0620",	x"0740",
	x"0380",	x"0380",	x"0380",	x"0380",	x"0380",	x"0fe0",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"3ffe",	x"301c",	x"2038",	x"0070",	x"00e0",	x"01c0",
	x"0380",	x"0700",	x"0e02",	x"1c06",	x"381c",	x"7ffc",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"07c0",	x"0400",	x"0400",	x"0400",	x"0400",	x"0400",	x"0400",
	x"0400",	x"0400",	x"0400",	x"0400",	x"0400",	x"0400",	x"0400",	x"07e0"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"2000",	x"1000",	x"0800",	x"0400",	x"0200",	x"0100",
	x"0080",	x"0040",	x"0020",	x"0010",	x"0008",	x"0004",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"03e0",	x"0020",	x"0020",	x"0020",	x"0020",	x"0020",	x"0020",
	x"0020",	x"0020",	x"0020",	x"0020",	x"0020",	x"0020",	x"0020",	x"07e0"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0fc0",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000"
),                                                                                            
                                                                                              
(                                                                                             
	                                                                                          
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"ffff",	x"0000"
),                                                                                            
                                                                                              
(	                                                                                          
	x"0000",	x"0000",	x"1800",	x"3000",	x"3800",	x"0000",	x"0000",	x"0000",
	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000"
),
   (
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"1ff0",	x"3818",--a
		x"0018",	x"0ff8",	x"3018",	x"6018",	x"707a",	x"1f9c",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"7800",	x"1800",	x"1800",	x"1800",	x"1ff8",	x"180e",
		x"1806",	x"1806",	x"1806",	x"1806",	x"1c0c",	x"13f0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0ffc",	x"301c",
		x"7000",	x"6000",	x"7000",	x"3002",	x"1c0c",	x"07f0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"00f8",	x"0018",	x"0018",	x"0018",	x"1ff8",	x"3018",
		x"6018",	x"6018",	x"6018",	x"6018",	x"3838",	x"0fde",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0ff8",	x"300c",
		x"300e",	x"7ff0",	x"7000",	x"3000",	x"1c0c",	x"03f0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"00f8",	x"0100",	x"0300",	x"0300",	x"0ff0",	x"0300",--f
		x"0300",	x"0300",	x"0300",	x"0300",	x"0300",	x"1fe0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"1fff",	x"3038",
		x"3018",	x"3038",	x"0ce0",	x"3300",	x"1fe0",	x"701c",	x"600e",	x"3ffc"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"f000",	x"3000",	x"3000",	x"3000",	x"37f8",	x"381c",
		x"301c",	x"301c",	x"301c",	x"301c",	x"301c",	x"fc3e",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0380",	x"0000",	x"0000",	x"0000",	x"0f80",	x"0180",
		x"0180",	x"0180",	x"0180",	x"0180",	x"0180",	x"0ff0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		X"0000",	X"0000",	X"0070",	X"0000",	X"0000",	X"0000",	X"01f0",	X"0070",--k
		X"0070",	x"0070",	X"0070",	X"0070",	X"0070",	X"0070",	X"0460",	X"07c0"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"7800",	x"1800",	x"1800",	x"1800",	x"1878",	x"1840",
		x"1980",	x"1fc0",	x"18e0",	x"1870",	x"1838",	x"7e7e",	x"0000",	x"0000"
	),                                                                                      
	(                                                          
		x"0000",	x"0000",	x"0f80",	x"0180",	x"0180",	x"0180",	x"0180",	x"0180",
		x"0180",	x"0180",	x"0180",	x"0180",	x"0180",	x"0ff0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"fffc",	x"718e",
		x"718e",	x"718e",	x"718e",	x"718e",	x"718e",	x"fbdf",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"7ff8",	x"3818",
		x"381c",	x"381c",	x"381c",	x"381c",	x"381c",	x"7c3e",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"1ff8",	x"300c",--p
		x"6006",	x"6006",	x"6006",	x"7006",	x"381c",	x"07e0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"7ff8",	x"180c",
		x"1806",	x"1806",	x"1806",	x"1806",	x"1c0c",	x"1bf0",	x"1800",	x"7f00"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"1ff8",	x"3018",
		x"6018",	x"6018",	x"6018",	x"7018",	x"3838",	x"0fd8",	x"0018",	x"007e"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"7cfe",	x"0f00",
		x"0c00",	x"0c00",	x"0c00",	x"0c00",	x"0c00",	x"7f80",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"1ffc",	x"1804",
		x"1e00",	x"07f0",	x"001c",	x"200e",	x"180c",	x"17f0",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0100",	x"0100",	x"0300",	x"1ff8",	x"0300",
		x"0300",	x"0300",	x"0300",	x"0300",	x"0384",	x"01f8",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"703c",	x"301c",
		x"301c",	x"301c",	x"301c",	x"301c",	x"383c",	x"0fde",	x"0000",	x"0000"
	),                                                                                       
	(                                                                                        
		X"0000",	X"0000",	X"0000",	X"0000",	X"0000",	X"0000",	X"781c",	X"1808",
		X"0c10",	X"0e20",	X"0620",	X"0340",	X"0380",	X"0180",	X"0000",	X"0000"
	),                                                                                      
	(                                                          
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"6186",	x"3184",
		x"31cc",	x"1bc8",	x"1a68",	x"1a70",	x"0c70",	x"0c30",	x"0000",	x"0000"
	),                                                                                        
	(                                                                                         
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"3c1c",	x"0e20",
		x"0340",	x"0180",	x"02c0",	x"0c70",	x"1018",	x"7c7e",	x"0000",	x"0000"
	),                                                                                        
	(                                                                                         
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"383c",	x"1810",
		x"0c20",	x"0e20",	x"0640",	x"0380",	x"0380",	x"0100",	x"0300",	x"7c00"
	),                                                                                        
	(                                                                                         
		x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"0000",	x"3ffc",	x"2038",--z
		x"00e0",	x"01c0",	x"0700",	x"0e04",	x"380c",	x"7ffc",	x"0000",	x"0000"
	)                                                                     
);
type oled_num_32x32 is array (0 to 9,0 to 31) of std_logic_vector(0 to 31);
constant num_table2:oled_num_32x32:=
(	
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"0007E000",X"001E7800",X"001C3800",--0
	X"003C3C00",X"00381C00",X"00381C00",X"00781E00",X"00781E00",X"00700E00",X"00700E00",X"00700E00",
	X"00700E00",X"00700E00",X"00700E00",X"00781E00",X"00781E00",X"00381C00",X"00381C00",X"003C3C00",
	X"001C3800",X"000E7000",X"0007E000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"0001C000",X"0007C000",X"001FC000",--1
	X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",
	X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",
	X"0003C000",X"0003C000",X"000FF800",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001DF000",X"00387800",--2
	X"00303800",X"00303C00",X"00703C00",X"00603C00",X"00003C00",X"00003800",X"00003800",X"00007800",
	X"00007000",X"0000E000",X"0000E000",X"0001C000",X"00038000",X"00070000",X"000E0000",X"000C0E00",
	X"001C0C00",X"003FFC00",X"007FFC00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001CF000",X"00387800",--3
	X"00303800",X"00303800",X"00003800",X"00003000",X"00007000",X"0000E000",X"0003E000",X"000FF800",
	X"00007800",X"00003C00",X"00001C00",X"00001C00",X"00001C00",X"00001C00",X"00001800",X"00003800",
	X"00003000",X"007CE000",X"003FC000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00007000",X"00007000",X"0000F000",--4
	X"0001F000",X"0001F000",X"0003F000",X"00037000",X"00077000",X"000E7000",X"000C7000",X"001C7000",
	X"00187000",X"00387000",X"00707000",X"00607000",X"007FFE00",X"00007000",X"00007000",X"00007000",
	X"00007000",X"00007000",X"00007000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000C00",X"0007FC00",X"0007F800",X"000E0000",--5
	X"000E0000",X"001C0000",X"001C0000",X"001F8000",X"003FC000",X"0037E000",X"0000F000",X"00007800",
	X"00003800",X"00003800",X"00001C00",X"00001C00",X"00001C00",X"00001800",X"00003800",X"00003800",
	X"00007000",X"007CE000",X"003FC000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000C00",X"0000FC00",X"0001C000",X"00078000",--6
	X"000F0000",X"000E0000",X"001E0000",X"001C0000",X"003C0000",X"003FF000",X"007E7800",X"00783C00",
	X"00781E00",X"00781E00",X"00701E00",X"00700E00",X"00780E00",X"00380E00",X"00380E00",X"00381C00",
	X"001C1C00",X"000E3800",X"0007F000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"003FFC00",X"003FFC00",X"00301C00",--7
	X"00701800",X"00603800",X"00003800",X"00003800",X"00003000",X"00007000",X"00007000",X"00007000",
	X"0000E000",X"0000E000",X"0000E000",X"0001C000",X"0001C000",X"0001C000",X"0003C000",X"00038000",
	X"00038000",X"00038000",X"00070000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FF000",X"001C3800",X"00381800",--8
	X"00381C00",X"00381C00",X"00381C00",X"003C3800",X"001C3800",X"001F7000",X"000FC000",X"0007E000",
	X"0007F000",X"000EF800",X"001C7800",X"00383C00",X"00381C00",X"00381C00",X"00381C00",X"00381C00",
	X"003C1C00",X"001C3800",X"000FF000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001C7000",X"00383800",--9
	X"00383C00",X"00781C00",X"00701C00",X"00701C00",X"00701E00",X"00781E00",X"00781E00",X"00381E00",
	X"003C1C00",X"001E7C00",X"000FFC00",X"00003C00",X"00003800",X"00007800",X"0000F000",X"0000E000",
	X"0001C000",X"00078000",X"003E0000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	)                                                                                  
);
type LCD_lux is array (0 to 2,0 to 31) of std_logic_vector(0 to 31);
constant lux_table:LCD_lux:=
(
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"01FF0000",X"00780000",X"00780000",
	X"00780000",X"00780000",X"00780000",X"00780000",X"00780000",X"00780000",X"00780000",X"00780000",
	X"00780000",X"00780000",X"00780000",X"00780000",X"00780000",X"00780380",X"00780300",X"00780700",
	X"00780F00",X"00783F00",X"01FFFE00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"07FC3FC0",X"01E00E00",X"01E00E00",
	X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",
	X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00E00",X"00E00C00",X"00F01C00",
	X"00701800",X"00783800",X"001FE000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"03FF3FC0",X"00F80F00",X"00780E00",
	X"003C0E00",X"001C1C00",X"001E3800",X"000E3000",X"000F7000",X"0007E000",X"0003C000",X"0003C000",
	X"0003E000",X"0007E000",X"0006F000",X"000E7000",X"001C7800",X"00183C00",X"00383C00",X"00701E00",
	X"00F01E00",X"01F01F00",X"07F87FE0",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	)
);
type LCD_colon is array (0 to 1,0 to 31) of std_logic_vector(0 to 31);
constant colon_table:LCD_colon:=
(
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
	X"0003C000",X"0003C000",X"0003C000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
	X"00000000",X"00000000",X"00000000",X"00000000",X"0003C000",X"0003C000",X"0003C000",X"00000000",
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	)
);
type LCD_tep is array (0 to 2,0 to 31) of std_logic_vector(0 to 31);
constant tep_table:LCD_tep:=
(
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"01FFFF00",X"01E38F00",X"01C38700",
	X"01838300",X"01838300",X"01038000",X"00038000",X"00038000",X"00038000",X"00038000",X"00038000",
	X"00038000",X"00038000",X"00038000",X"00038000",X"00038000",X"00038000",X"00038000",X"00038000",
	X"00038000",X"0007C000",X"001FF000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"01FFFE00",X"00781E00",X"00780E00",
	X"00780600",X"00780600",X"00780000",X"00780000",X"00781800",X"00781800",X"00783800",X"007FF800",
	X"00783800",X"00781800",X"00781800",X"00780000",X"00780000",X"00780000",X"00780380",X"00780700",
	X"00780700",X"00781F00",X"01FFFE00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00FFE000",X"003C7C00",X"003C1E00",
	X"003C0E00",X"003C0F00",X"003C0F00",X"003C0F00",X"003C0F00",X"003C0F00",X"003C1E00",X"003C3C00",
	X"003FF800",X"003C0000",X"003C0000",X"003C0000",X"003C0000",X"003C0000",X"003C0000",X"003C0000",
	X"003C0000",X"003E0000",X"00FF8000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	)
);
type oled_num2_32x32 is array (0 to 10,0 to 31) of std_logic_vector(0 to 31);
constant num_table3:oled_num2_32x32:=
(	
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"0007E000",X"001E7800",X"001C3800",--0
	X"003C3C00",X"00381C00",X"00381C00",X"00781E00",X"00781E00",X"00700E00",X"00700E00",X"00700E00",
	X"00700E00",X"00700E00",X"00700E00",X"00781E00",X"00781E00",X"00381C00",X"00381C00",X"003C3C00",
	X"001C3800",X"000E7000",X"0007E000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"0001C000",X"0007C000",X"001FC000",--1
	X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",
	X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",X"0001C000",
	X"0003C000",X"0003C000",X"000FF800",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001DF000",X"00387800",--2
	X"00303800",X"00303C00",X"00703C00",X"00603C00",X"00003C00",X"00003800",X"00003800",X"00007800",
	X"00007000",X"0000E000",X"0000E000",X"0001C000",X"00038000",X"00070000",X"000E0000",X"000C0E00",
	X"001C0C00",X"003FFC00",X"007FFC00",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001CF000",X"00387800",--3
	X"00303800",X"00303800",X"00003800",X"00003000",X"00007000",X"0000E000",X"0003E000",X"000FF800",
	X"00007800",X"00003C00",X"00001C00",X"00001C00",X"00001C00",X"00001C00",X"00001800",X"00003800",
	X"00003000",X"007CE000",X"003FC000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"00007000",X"00007000",X"0000F000",--4
	X"0001F000",X"0001F000",X"0003F000",X"00037000",X"00077000",X"000E7000",X"000C7000",X"001C7000",
	X"00187000",X"00387000",X"00707000",X"00607000",X"007FFE00",X"00007000",X"00007000",X"00007000",
	X"00007000",X"00007000",X"00007000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000C00",X"0007FC00",X"0007F800",X"000E0000",--5
	X"000E0000",X"001C0000",X"001C0000",X"001F8000",X"003FC000",X"0037E000",X"0000F000",X"00007800",
	X"00003800",X"00003800",X"00001C00",X"00001C00",X"00001C00",X"00001800",X"00003800",X"00003800",
	X"00007000",X"007CE000",X"003FC000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000C00",X"0000FC00",X"0001C000",X"00078000",--6
	X"000F0000",X"000E0000",X"001E0000",X"001C0000",X"003C0000",X"003FF000",X"007E7800",X"00783C00",
	X"00781E00",X"00781E00",X"00701E00",X"00700E00",X"00780E00",X"00380E00",X"00380E00",X"00381C00",
	X"001C1C00",X"000E3800",X"0007F000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"003FFC00",X"003FFC00",X"00301C00",--7
	X"00701800",X"00603800",X"00003800",X"00003800",X"00003000",X"00007000",X"00007000",X"00007000",
	X"0000E000",X"0000E000",X"0000E000",X"0001C000",X"0001C000",X"0001C000",X"0003C000",X"00038000",
	X"00038000",X"00038000",X"00070000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                   
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FF000",X"001C3800",X"00381800",--8
	X"00381C00",X"00381C00",X"00381C00",X"003C3800",X"001C3800",X"001F7000",X"000FC000",X"0007E000",
	X"0007F000",X"000EF800",X"001C7800",X"00383C00",X"00381C00",X"00381C00",X"00381C00",X"00381C00",
	X"003C1C00",X"001C3800",X"000FF000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),                                                                                            
	(                                                                                             
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"000FE000",X"001C7000",X"00383800",--9
	X"00383C00",X"00781C00",X"00701C00",X"00701C00",X"00701E00",X"00781E00",X"00781E00",X"00381E00",
	X"003C1C00",X"001E7C00",X"000FFC00",X"00003C00",X"00003800",X"00007800",X"0000F000",X"0000E000",
	X"0001C000",X"00078000",X"003E0000",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	),
	(
	X"00000000",X"00000000",X"00000000",X"00000000",X"00000000",X"03FE7FC0",X"00F00F00",X"00700F00",--H
	X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"007FFF00",
	X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",X"00700F00",
	X"00F00F00",X"00F81F00",X"03FE7FC0",X"00000000",X"00000000",X"00000000",X"00000000",X"00000000"
	)
);
type oled_pic_16x16 is array (0 to 1,0 to 15) of std_logic_vector(0 to 15);
constant pic_table3:oled_pic_16x16:=
(
	(
	   X"0000",	X"07e0",	X"0ff0",	X"1818",	X"380c",	X"300c",	X"6006",	X"6006",   --�f��
	   X"6006",	X"6006",	X"300c",	X"300c",	X"1918",	X"0f30",	X"0700",	X"0f00"	   
	),
	(
	   X"0000",	X"07e0",	X"0ff0",	X"1818",	X"380c",	X"300c",	X"6006",	X"6006",   --����
	   X"6006",	X"6006",	X"300c",	X"300c",	X"1898",	X"0cf0",	X"00e0",	X"00f0"		   
	)
);
------------------------------------------------------------------------TSL2561
SIGNAL  TSL2561_data : STD_LOGIC_VECTOR(14 DOWNTO 0);
SIGNAL  TSL2561_int  :integer range 0 to 9999;            
SIGNAL  d0, d0_last  :integer range 0 to 9999;   
SIGNAL  lx1,lx2,lx3,lx4,lx5 :integer range 0 to 9;   	                                
------------------------------------------------------------------------------------------DHT11
SIGNAL HU_BUFF, TE_BUFF : STD_LOGIC_VECTOR(7 DOWNTO 0); 
signal TE,HU:integer range 0 to 255; 
SIGNAL DHT11_error : STD_LOGIC;   
---------------------------------------------------------------------------------------------------KEYBOARD
--SIGNAL keyin,keyin_last : std_logic_vector(0 to 15);
signal pb:std_logic_vector(3 downto 0);
signal pe,per:std_logic;
signal swr:std_logic_vector(7 downto 0);

SIGNAL event_S1, event_S2, event_S3, event_S4, event_S5 , event_S6: STD_LOGIC;        
---------------------------------------------------------------------------------------------------7SEG
signal seg1:std_logic_vector(3 downto 0);
signal seg2:std_logic_vector(3 downto 0);
signal c1015:std_logic_vector(7 downto 0);
type seg_ram is array(0 to 7)of integer range 0 to 15;
signal segr :seg_ram;
type seg_rom is array(0 to 15)of std_logic_vector(6 downto 0);
signal seg_num :seg_rom:=
(
	"1111110" ,"0110000" ,"1101101" ,"1111001" ,"0110011" ,"1011011" ,"0011111" ,"1110000" 
	,"1111111" ,"1110011" ,"1110111" ,"0011111" ,"1001110" ,"0111101" ,"1001111" ,"0000000"
);
------------------------------------------------------------------------------------dot8*8
type dot_type is array (0 to 7) of std_logic_vector(7 downto 0);
signal dotR : dot_type;
signal dotG : dot_type;
signal coml : dot_type:=(X"80",X"40",X"20",X"10",X"08",X"04",X"02",X"01");
type code is array (0 to 15) of std_logic_vector(63 downto 0);
signal num : code:=(
"0000000000011000001001000010010000100100001001000001100000000000",--0
"0000000000001000000110000000100000001000000010000000100000000000",--1
"0000000000011000001001000000010000001000000100000011110000000000",--2
"0000000000011000001001000000010000011000000001000010010000011000",--3
"0000000000001000000110000010100000101000001111000000100000000000",--4
"0000000000111100001000000011100000000100000001000011100000000000",--5
"0000000000011000001000000011100000100100001001000001100000000000",--6
"0000000000111100001001000000010000001000000010000000100000000000",--7
"0000000000011000001001000010010000111100001001000010010000011000",--8
"0000000000011000001001000010010000011100000001000010010000011000",--9
x"001824243c242400", --A
x"0038243824380000", --B
x"0018204040201800", --C
x"0030282424283000", --D
x"0078407840407800", --E
x"0078407840404000"  --F
);
--------------------------------------------------------------------------------------------------SD178B  
--SIGNAL  sd178_ena, sd178_rw, sd178_busy, sd178_ack_error  : std_logic;   
--SIGNAL  sd178_addr      : STD_LOGIC_VECTOR(6 DOWNTO 0);     
--SIGNAL  cnt_byte   :integer range 0 to 30; 
--SIGNAL  var_vol,var_vol_last  :integer range 0 to 9; 
signal sd178_ena, sd178_rw, sd178_busy : std_logic;
signal sd178_data_wr, sd178_data_rd : std_logic_vector(7 downto 0);
signal sdbyte : integer range 0 to 31;	--�X�r��
signal sdtime,sdtimer: std_logic;				--����
signal sdsub : integer range 0 to 3;	--SD����
signal sd_t : integer range 0 to 15_000_000;
signal sdmode: integer range 0 to 10;
signal sound:std_logic_vector(7 downto 0);
signal sd_speed:std_logic_vector(7 downto 0);
signal channel:integer range 0 to 3;
signal srun,srunr:std_logic;
signal remode:integer range 0 to 5;
type word_ram is array(0 to 19)of std_logic_vector(7 downto 0);                                
signal word_buf : word_ram:=( x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
--x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
 --"�ЧA���n����" x"BD",x"D0",x"A7",x"41",x"B0",x"B5",x"A6",x"6E",x"C1",x"C2",x"C1",x"C2",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
 --rt x"B7",x"4F",x"B7",x"4F",x"AD",x"44",x"AD",x"44",x"AF",x"75",x"A5",x"69",x"B7",x"52",x"BC",x"4B",x"BC",x"4B",x"00",x"00");
type wordnum_rom is array(0 to 9,0 to 1)of std_logic_vector(7 downto 0);
signal wordnum : wordnum_rom :=(
	( x"B9",x"73"),	( x"A4",x"40"),	( x"A4",x"47"),	( x"A4",x"54"),( x"A5",x"7C"),( x"A4",x"AD"),( x"A4",x"BB"),	
	
	( x"A4",x"43"),( x"A4",x"4B"),( x"A4",x"45")
);


-------------------------------------------------------------------------------------------other
--ck signal
signal q : std_logic_vector(25 downto 0);
signal ck_1M 	: std_logic;
signal ck_LCD 	: std_logic;
signal ck_b		: std_logic;
signal ck_pb	: std_logic;
signal bp		: std_logic_vector(1 downto 0);
signal ck_bz	: std_logic;
signal ck_mot	:std_logic;
signal ck_1s	:std_logic;
---------------------------------------
signal rst:std_logic;
---------------------------------------------------------------       
SIGNAL  d3 :integer range 0 to 20; 

-------------------------------------------------------------------------------------------motor
SIGNAL  mode_motor :integer range 0 to 10;
SIGNAL  motor_speed1,motor_speed2   :integer range 0 to 10;
SIGNAL  motor_dir1,motor_dir2 : STD_LOGIC;   --�����౱��     
-------------------------------------------------------------------------------------------LCD   
SIGNAL  clk: STD_LOGIC;
SIGNAL  x  :integer range 0 to 127; 
SIGNAL  y  :integer range 0 to 255; 
SIGNAL  d  :integer range 0 to 15;      
SIGNAL  fsm,fsm_back,fsm_back2   :integer range 0 to 150;
SIGNAL  address: STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL  RGB : STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL  add : STD_LOGIC_VECTOR(14 DOWNTO 0);
SIGNAL  e : STD_LOGIC_VECTOR(2 DOWNTO 0);
SIGNAL  data_out ,RGB_data,LCD_t  : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL  DC_data    : std_logic;   
-------------------------------------------------------------------------------------------RAM
SIGNAL we2   : std_logic;
SIGNAL a2     : std_logic_vector(14 downto 0);
SIGNAL di2, do2 : std_logic_vector(5 downto 0);
-------------------------------------------------------------------------------------------RS
Type mem is array(0 to 1)of std_logic_vector(7 downto 0);
signal dataR : mem;
Type mFm is array(0 to 7)of std_logic_vector(7 downto 0);--32byte
signal dataT : mfm;


signal 	PcOkFlag ,flag ,bt,btt : std_logic;
--===============================================================�{��
signal seg_a,seg_s:std_logic;

--Type password is array(0 to 5,0 to 3)of std_logic_vector(3 downto 0);
--signal pass,ans,passspace : password:=
--(
--	(x"0", x"0", x"0", x"0"),(x"0", x"0", x"0", x"0"),
--	(x"0", x"0", x"0", x"0"),(x"0", x"0", x"0", x"0"),
--	(x"0", x"0", x"0", x"0"),(x"0", x"0", x"0", x"0")
--);
--
--Type timeram is array(0 to 5)of integer range 0 to 9999;
--signal secram : timeram;


--signal 
--=========================================
begin  



main:process(ck)            
variable t,ts,tt,ttt,sdt:integer range 0 to 15_000_000;
variable start,startr:std_logic;
----------------------------------------------
variable LD: integer range 0 to 10;--std_logic_vector(3 downto 0); --
variable lx1r,lx2r,lx3r,lx4r,lx5r: integer range 0 to 9;
----------------------------------------------
variable tr1,tr2,tr3,tr4,tr5: integer range 0 to 37;
----------------------------------------------
variable R,G,B:std_logic_vector(4 downto 0);
--variable remain :integer range 0 to 4:=4;
--variable remain1,remain2,remain3,remain4 :integer range 0 to 1;
variable op,c:integer range 0 to 10;
variable LEDH:integer range 0 to 6;
-------------------------------------------
variable choose:integer range 0 to 3;
variable vol,spd:integer range 0 to 5;
-------------------------------------
variable color:integer range 0 to 10;
variable colorR,colorG,colorB:integer range 0 to 3;
variable mode:integer range 0 to 3;
variable ks:integer range 0 to 3;
variable j:integer range 0 to 160;
variable first:integer range 0 to 1;
variable Rs:integer range 0 to 3;

begin
--
--if rising_edge(ck_1s) then
--	
--end if;


if rising_edge(ck_1M) then
per<=pe;
--bt<='0';
--seg_s<='1';
LED<=not x"0000";

if per='0' and pe='1' then
	if pb=0 then
		c:=1;
		t:=0;
		start:='1';
	end if;
	if pb=2 then
		c:=0;
		start:='0';
		t:=0;
	end if;
end if;

			
segr<=(TE/10, TE mod 10, 0, 12, conv_integer(motor_speed1)/10, conv_integer(motor_speed1)mod 10, 0, 0);

--motor_speed1<=5;
--motor_dir1<='0';
--for i in 0 to 7 loop
--	dotR(i)<=num(0)((i+1)*8-1 downto i*8);
--	dotG(i)<=num(1)((i+1)*8-1 downto i*8);
--end loop;

if swr/=sw then
	swr<=sw;
	c:=0;t:=0;
else
case t is
when 0=>--t:=1_000_000;
--------------------------------------------------------
	case c is
		when 0=>rst<='0';	--reset
				seg_s<='0';
				LD:=0;
				motor_speed1<=0;
				start:='0';
				
				choose:=0;
				vol:=3;spd:=0;
				c:=10;
				
				color:=0;colorR:=0;colorG:=0;colorB:=0;
				ks:=0;
				first:=0;
				RS:=0;
				
		when 1=> 	--start?
					case swr(7 downto 6) is
						when "00"=>c:=2;	LD:=0;
						when "01"=>c:=3;	LD:=1;seg_s<='1';TE<=conv_integer(TE_buff);
						when "10"=>c:=4;	LD:=1;
						when "11"=>c:=5;	
					end case;
				
		when 2=>if start='1' then
					t:=500_000;
					case color is
						when 0=>color:=1;LD:=1;
						when 1=>LD:=0;
								if ks<2 then
									ks:=ks+1;
									color:=0;
								else
									ks:=0;
									color:=2;
								end if;
						when 2=>t:=2_000_000;
								color:=0;LD:=2;
						when others=>null;
					end case;
				end if;
		when 3=>if start='1' then
					if first=0 then
						first:=1;
						motor_speed1<=3;
					end if;
					if TE/=te_buff then
						if TE>TE_buff then
							motor_speed1<=motor_speed1-1;
						else
							motor_speed1<=motor_speed1+1;
						end if;
						TE<=conv_integer(TE_buff);
					end if;
					LD:=3;
					if j<160 then
						j:=j+1;
					else
						j:=0;
					end if;
					t:=50_000;
				else
					motor_speed1<=0;first:=0;
				end if;
		when 4=>if start='1' then
					t:=1_000_000;
					lx2r:=lx2;lx3r:=lx3;lx4r:=lx4;lx5r:=lx5;
					LD:=4;
					if TSL2561_int<20 then
						motor_dir1<='1';
						if RS>0 then Rs:=Rs-1; else Rs:=3; end if;
					else
						motor_dir1<='0';
						if RS<3 then Rs:=Rs+1; else Rs:=0; end if;
					end if;
					motor_speed1<=5;
				else
					motor_speed1<=0;
				end if;
		when 5=>if start='1' then
					LD:=5;
					if sdmode=10 then
						sdmode<=1;
					end if;
					if per='0' and pe='1' then
						if pb=4 then
							case choose is
								when 1=>if vol<5 then vol:=vol+1; end if;
								when 2=>if spd<5 then spd:=spd+1; end if;
								when 3=>if channel<2 then channel<=channel +1; else channel<=0; end if;
								when others=>null;
							end case;
						end if;
						if pb=5 then
							case choose is
								when 1=>if vol>0 then vol:=vol-1; end if;
								when 2=>if spd>0 then spd:=spd-1; end if;
								when 3=>if channel>0 then channel<=channel -1; else channel<=2; end if;
								when others=>null;
							end case;
						end if;
						if pb=6 then
							sdt:=1;
							sd_t<=0;
							sdsub<=0;
							remode<=1;
							sdmode<=0;
							sound<=conv_std_logic_vector((159 + vol*10),8);
							sd_speed<=conv_std_logic_vector((spd*5),8);
						end if;
						if pb=12 then
							choose:=choose+1;
						end if;

					end if;

				end if;
		when others=>null;
	end case;
		
--------------------------------------------------------		
when others=>t:=t-1;
end case;
end if;
--case ts is
--	when 0=>case LEDH is
--				when 0=>LED_R<='0';
--						LED_G<='0';
--						LED_Y<='0';
--						LED_RGB<="000";
--						--ts:=1_000_000;LEDH:=LEDH+1;
--				
--				when others=>null;
--			end case;
--	when others=>ts:=ts-1;
--end case;

case LD is	
	when 0=>RGB<="0000000000000000";
	when 1=>RGB<="1111111111111111";

	when 2=>RGB<=conv_std_logic_vector(x/4,5)& conv_std_logic_vector(y/5,5)&"000000";
		
			---------------------------------------------------------------------
--			elsif (y>=26*1 and y<26*2) or (y>=26*3 and y<26*4) or (y>=26*5 and y<26*6) then
--					if (y>=26*id and y<26*(id+1)) then
--						if (x>0 and x<jk) then
--							RGB<="0000000000011111";
--						else
--							RGB<="0000001010000000";
--						end if;
--					else
--						RGB<="0000011111000000";
--					end if;
--							
--			else
--				RGB<="0000000000000000";
--			end if;
	when 3=>if j<160-32 then
				if (y>j and y<=j+32) then
					if (((x>32*0 and x<=32*1) and num_table2(TE/10,y-j)(x-32*0)='1') or
						((x>32*1 and x<=32*2) and num_table2(TE mod 10,y-j)(x-32*1)='1') 
					) then                                  
						RGB<="0000001111100000";
					else
						RGB<="1111111111111111";
					end if;
				end if;
			else
				if (y>j or y<=j+32-160) then
					if y>j then
						if (((x>32*0 and x<=32*1) and num_table2(TE/10,y-j)(x-32*0)='1') or
							((x>32*1 and x<=32*2) and num_table2(TE mod 10,y-j)(x-32*1)='1') 
						) then                                  
							RGB<="0000001111100000";
						else
							RGB<="1111111111111111";
						end if;
					else
						if (((x>32*0 and x<=32*1) and num_table2(TE/10,y-j)(x-32*0)='1') or
							((x>32*1 and x<=32*2) and num_table2(TE mod 10,y-(j))(x-32*1)='1') 
						) then                                  
							RGB<="0000001111100000";
						else
							RGB<="1111111111111111";
						end if;
					end if;
				end if;
			end if;
	when 4=>if (y>32*0 and y<=32*1) then
				if (((x>32*0 and x<=32*1) and num_table2(lx2r,y-32*0)(x-32*0)='1') or
					((x>32*1 and x<=32*2) and num_table2(lx3r,y-32*0)(x-32*1)='1') or
					((x>32*2 and x<=32*3) and num_table2(lx4r,y-32*0)(x-32*2)='1') or
					((x>32*3 and x<=32*3+2) and (y>30 and y<=32)) or
					((x>32*3 and x<=32*4) and num_table2(lx5r,y-32*0)(x-32*3)='1')
				) then                                  
					if (lx2r*1000+lx3r*100+lx4r*10+lx5r)<20 then
						RGB<="0000001111100000";
					else
						RGB<="0000000000000000";
					end if;
				else
					RGB<="1111111111111111";
				end if;
			elsif (y>32*1 and y<=16*3) then
				case Rs is
					when 0=>if (((x>16*0 and x<=16*1) and num_table1(82,y)(x)='1')) then
								RGB<="0000000000000000";
							else
								RGB<="1111111111111111";
							end if;
					when 1=>if (((x>16*0 and x<=16*1) and num_table1(82,x)(16-y)='1')) then
								RGB<="0000000000000000";
							else
								RGB<="1111111111111111";
							end if;
					when 2=>if (((x>16*0 and x<=16*1) and num_table1(82,16-y)(16-x)='1')) then
								RGB<="0000000000000000";
							else
								RGB<="1111111111111111";
							end if;
					when 3=>if (((x>16*0 and x<=16*1) and num_table1(82,16-x)(y)='1')) then
								RGB<="0000000000000000";
							else
								RGB<="1111111111111111";
							end if;
				end case;
			else
				RGB<="1111111111111111";	
			end if;
	when 5=>if (y>0 and y<=50) then
				if (((y>16*0 and y<=16*1) and (x>16*0 and x<=16*1) and num_table1(86,y-16*0)(x-16*1)='1') or--
					((y>16*0 and y<=16*1) and (x>16*1 and x<=16*2) and num_table1(111,y-16*0)(x-16*2)='1') or
					((y>16*0 and y<=16*1) and (x>16*2 and x<=16*3) and num_table1(108,y-16*0)(x-16*3)='1') or
					((y>16*0 and y<=16*1) and (x>16*3 and x<=16*4) and num_table1(58,y-16*0)(x-16*4)='1') or
					((y>16*0 and y<=16*1) and (x>16*4 and x<=16*5) and num_table1(vol+48,y-16*0)(x-16*5)='1') 
				) then             
					RGB<="0000000000000000";
				else
					if choose=1 then
						RGB<="1011100000000000";
					else
						RGB<="1111100000000000";
					end if;
				end if;
			elsif (y>50 and y<=100) then
				if (((y>50 and y<=50+16) and (x>16*0 and x<=16*1) and num_table1(115,y-50)(x-16*1)='1') or--
					((y>50 and y<=50+16) and (x>16*1 and x<=16*2) and num_table1(112,y-50)(x-16*2)='1') or
					((y>50 and y<=50+16) and (x>16*2 and x<=16*3) and num_table1(100,y-50)(x-16*3)='1') or
					((y>50 and y<=50+16) and (x>16*3 and x<=16*4) and num_table1(58 ,y-50)(x-16*4)='1') or
					((y>50 and y<=50+16) and (x>16*4 and x<=16*5) and num_table1(spd+48,y-50)(x-16*5)='1') 
				) then             
					RGB<="0000000000000000";
				else
					if choose=2 then
						RGB<="0000010111000000";
					else
						RGB<="0000011111000000";
					end if;
				end if;
			else
				if choose=3 then
					RGB<="0000000000010111";
				else
					RGB<="0000000000011111";
				end if;
				
				
				if channel <2 then
					if (((y>100 and y<=116) and (x>16*0 and x<=16*1) and num_table1(82,y-100)(x-16*0)='1') )
					then
						RGB<="0000000000000000";
					end if;
				end if;	
				if channel/=1 then
					if (((y>100 and y<=116) and (x>16*1 and x<=16*2) and num_table1(76,y-100)(x-16*1)='1') )
					then
						RGB<="0000000000000000";
					end if;
				end if;		
					
				
					
				--end if;
			end if;
	when others=>null;		
end case;
		
----------------------------------------------------------------------	
if rst='0' then
rst<='1';
sdt:=1;
sd_t<=0;
sdsub<=0;
sdtime<='0';
remode<=0;
sdmode<=0;
sound<=x"C2";
channel<=0;
sd_speed<=x"00";
else
case sdt is
when 0=>
----------------------------------------------------------------------
case sdsub is
	when 0=>
----------------------------------------------------------------------			
	case remode is
		when 0=>word_buf(0 to 1)<=(x"80",x"00");--reset
				sdbyte<=2;
				sdsub<=1;
				sd_t<=100_000;
				remode<=1;
		when 1=>LED_RGB<=LED_RGB+1;
			case channel is
				when 0=>word_buf(0 to 1)<=(x"8B", x"08");--���n�D07
						sdbyte<=2;
						sdsub<=1;
						sd_t<=50_000;
				when 1=>word_buf(0 to 1)<=(x"8B", x"0A");--�k�n�D06
						sdbyte<=2;
						sdsub<=1;
						sd_t<=50_000;
				when 2=>word_buf(0 to 1)<=(x"8B", x"09");--���n�D05
						sdbyte<=2;
						sdsub<=1;
						sd_t<=50_000;
				when others=>null;
--				when 3=>word_buf(0 to 1)<=(x"8B", x"01");--�L�n�D01
--						sdbyte<=2;
--						sdsub<=1;
--						sd_t<=50_000;
			end case;		

			remode<=2;
		
		when 2=>
			word_buf(0 to 1)<=(x"86" ,sound);--���q
			sdbyte<=2;
			sdsub<=1;
			sd_t<=50_000;
			remode<=3;
		when 3=>
			word_buf(0 to 1)<=(x"83" ,sd_speed);--�t��
			sdbyte<=2;
			sdsub<=1;
			sd_t<=50_000;
			remode<=4;
		when 4=>
			
			word_buf(0 to 1)<=(x"8F" ,"0000000" & start);--stop
			sdbyte<=2;
			sdsub<=1;
			sd_t<=100_000;
			
			remode<=5;
		when 5=>
			if startr/=start then
				startr:=start;
				remode<=4;
			else
			
----------------------------------------------------------
	case sdmode is
		when 0=>
				word_buf(0 to 1)<=(x"80",x"00");--reset
				sdbyte<=2;
				sdsub<=1;
				sd_t<=100_000;
				sdmode<=10;
				
		when 1=>word_buf(0 to 19)<=(x"A8", x"74", x"B2", x"CE", x"B6", x"7D", x"BE", x"F7",x"BC", x"B7", x"A9", x"F1",wordnum(conv_integer(TE_buff)/10,0),wordnum(conv_integer(TE_buff)/10,1),wordnum(conv_integer(TE_buff)mod 10,0),wordnum(conv_integer(TE_buff)mod 10,1),x"AB", x"D7", x"43",x"00");
				sdbyte<=20;
				sdsub<=1;
				sd_t<=7_000_000;
				
				sdmode<=3;
--		when 2=>word_buf(0 to 11)<=(
--				
--				sdbyte<=12;
--				sdsub<=1;
--				sd_t<=4_000_000;
--				
--				sdmode<=3;
		when 3=>word_buf(0 to 1)<=(wordnum(lx2,0),wordnum(lx2,1));
				word_buf(2 to 3)<=(wordnum(lx3,0),wordnum(lx3,1));
				word_buf(4 to 5)<=(wordnum(lx4,0),wordnum(lx4,1));
				word_buf(6 to 7)<=(x"C2", x"49");
				word_buf(8 to 9)<=(wordnum(lx5,0),wordnum(lx5,1));
				word_buf(10 to 15)<=(x"B0", x"C7", x"A7", x"4A", x"B4", x"B5");
				sdbyte<=16;
				sdsub<=1;
				sd_t<=3_000_000;
				
				sdmode<=4;
		when 4=>word_buf(0 to 4)<=(x"88", x"27", x"0E", x"00", x"01");
				sdbyte<=5;
				sdsub<=1;
				sd_t<=13_000_000;
				
				sdmode<=1;
		when others=>null;
	end case;
-----------------------------------------------------------------
			end if;
	end case;
-----------------------------------------------------
	when 1=>sdtime<='1';
			sdt:=200_000;
			sdsub<=2;
	when 2=>sdtime<='0';
			sdt:=sd_t;
			sdsub<=0;
			sd_t<=0;
	when others=>null;
end case;
-------------------------------------------------------------------------
when others=>sdt:=sdt-1;
end case;
end if;	
-------------------------------------------------------------------------		
end if;
      			
	   
end process;
-------------------------------------------------------------------------------------ck_maker
ck_macker:process(ck)
variable delay_100 : integer range 0 to 250_000;
variable delay_1s : integer range 0 to 25_000_000;
variable j : std_logic_vector(9 downto 0);
variable delay_1M : integer range 0 to 31;
begin

	if rising_edge(ck)then
		q <= q + 1;--ck maker

		if delay_1M = 25 then
			delay_1M := 0;
			ck_1M <= not ck_1M;
		else
			delay_1M := delay_1M + 1;
		end if;
		
		if delay_100 = 249_999 then
			delay_100 := 0;
			ck_mot <= not ck_mot;
		else
			delay_100 := delay_100 + 1;
		end if;
		
		if delay_1s = 24_999_999 then
			delay_1s := 0;
			ck_1s <= not ck_1s;
		else
			delay_1s := delay_1s + 1;
		end if;
		ck_LCD 	<= q(0);
		ck_b	<= q(19);
		ck_pb <=q(16);
		ck_bz <=q(17);
		
		--------------------------
		if j = "1111111111" then
			j := "0000000000";
		else
			j := not j(0) & j(9 downto 1);
		end if;
		
	end if;
-- 0 25M		-- 1 12.5M		-- 2 6.25M		-- 3 3.125M
-- 4 1.5625M	-- 5 781K		-- 6 390K		-- 7 195K
-- 8 97K		-- 9 48K		-- 10 24K		-- 11 12K
-- 12 6K		-- 13 3K		-- 14 1.5K		-- 15 762
-- 16 381		-- 17 190		-- 18 95		-- 19 47
-- 20 23		-- 21 11		-- 22 6			-- 23 3
-- 24 1.5		-- 25 0.7

end process;
--=================================================================================8*8
dot8x8:process(ck_1M)
variable c: integer range 0 to 7;
--variable RorG:std_logic;
begin

if rising_edge(ck_1M) then
	com<=coml(c);
	
--	case RorG is
--		when '0'=>
--		when '1'=>
--	end case;
	out_R<=not(dotR(c));
	out_G<=not(dotG(c));
	
	if c=7 then
		c:=0;
		--RorG:=not RorG;
	else
		c:=c+1;
	end if;
end if;
end process;
--==============================================================================
tsl:process(ck_1M)
variable cnt_step:integer range 0 to 1;
begin
if rising_edge(ck_1M) then
	case cnt_step is                                 --�ഫTSL2561��� 
		when 0=>TSL2561_int  <= CONV_INTEGER(TSL2561_data) mod 10000;
				cnt_step := 1;
		when 1=>cnt_step:=0;
				lx1 <= (TSL2561_int / 10000) mod 10;
				lx2 <= (TSL2561_int / 1000) mod 10;
				lx3 <= (TSL2561_int / 100) mod 10;
				lx4 <= (TSL2561_int / 10) mod 10;
				lx5 <= TSL2561_int mod 10;
	end case;
end if;
end process;
--==============================================================================
sd178_dri: process(ck)  --sd178
variable t      :integer range 0 to 50_000_000;       
variable cnt_loop       :integer range 0 to 50;       
variable cnt2,s178           :integer range 0 to 20;      
variable cnt_byte : integer range 0 to 31;
begin  
      if rising_edge(ck) then  --(ck'EVENT AND ck='1')  
		sdtimer<=sdtime;
		
         if(nReset='0')then 
            SD178_nrst <= '0'; 
            sd178_ena  <= '0';                                      
            s178   := 0;

         else
			if t=0 then
            CASE s178 IS  
               when 0=>  
                        SD178_nrst <= '1';
                        s178 := 1; 
 						t :=  12_000_000 ;           	--0.24��
               when 1=>  
                  
						--if (sdflag = '1') then 
						if (sdtime = '1' and sdtimer='0') then 
							cnt_byte := sdbyte;-- 18;           	           
							-- word_buf <= word2;     
							--word_buf <= w_1;  		
                            s178 :=2; 
                           -- led(15 downto 12) <= led(15 downto 12) + 1;
                        end if; 
                        --end if;
			   
               WHEN 2 =>                   
                                                
                        cnt2 := 0;
                        cnt_loop := 0;
                        s178 := 3;                                                                                                                               
                                                                       
               WHEN 3=>                                       --start write data

--                      sd178_addr      <= "0100000";               --write sd178_address 0x20
                        sd178_data_wr   <= word_buf(cnt_loop);	           --�󴫸��                         
                        sd178_rw        <= '0';                     --0/write  
                        s178      := 4;
                        
                        cnt_loop := cnt_loop + 1;                   --�ǰe��ƤW��+1 
               WHEN 4=>                      
                        sd178_ena   <= '1';                                                                    
                        s178  := 5;  

               WHEN 5=>                      
                        if sd178_busy = '1' then  
                            if cnt_loop >= cnt_byte  then 
                               sd178_ena    <= '0';
                               s178   := 7;                                                          
                            else                            
                               sd178_data_wr <= word_buf(cnt_loop);         --command    
                               sd178_rw      <= '0';                 --0/write                                                                                                                                                                             
                               cnt_loop := cnt_loop + 1;             --�ǰe��ƤW��+1
                               s178    := 6;
                           end if; 
                        end if;                         
               WHEN 6=>            
                        if sd178_busy = '0' then                             
                           sd178_ena    <= '0';                                                                                       
                           if cnt_loop >= cnt_byte  then                --cnt_byte �ǰe�ƶq
                              s178  := 7;   
                           else                           
                              s178    := 8;                                                                                                                                                                                                                                           
                           end if;          
                        end if; 
                           
               WHEN 8=>   s178 := 3;t:=500_000;     --delay10ms&redo
                           
               WHEN 7=>   s178 := 9;t:=10_000_000;   --delay0.2s&end

               WHEN 9=>                                   
						if (sdtime = '0') then                       
                            s178 :=0;
						end if;     
              when others =>                                          
                        s178    := 0;
                          
            END CASE;
         else t:=t-1;                  
		end if;
       end if;
      end if;    
end process;
--==============================================================================
key:process(ck_1M)
variable x: std_logic_vector(1 downto 0);
begin

if rising_edge(ck_pb) then
	case x is
		when "00"=> if ki/="1111"  then x:="01"; pb<="0000"; ko<="1110"; end if;
		when "01"=> if ki="1111" then ko<=ko(2 downto 0)& ko(3); pb<=pb+1;
					else x:="10"; pe<='1';
						if ki(3)<='0' then pb(3 downto 2)<="11";
						else pb(3 downto 2)<=not ki(2 downto 1);
						end if;  
					end if;
		when others=>if ki="1111" then x:="00"; ko<="0000";pe<='0'; end if; 
	end case;
end if;
end process;
--=================================================================
SEG_driver:process(ck)--�C�q��ܾ�
variable w:	integer range 0 to 7;
begin

if rising_edge(ck_1M) then

if seg_s='0' then
	segout_2<="00000000";
	segout	<="00000000";
else
	w:=w+1;
	if w>3 then
		seg1<=conv_std_logic_vector(segr(w),4);
	else
		seg2<=conv_std_logic_vector(segr(w),4);
	end if;
	
	if c1015=x"00" then
		seg_scan<=not x"01";
		c1015<=x"02";
	else
		c1015<= c1015(6 downto 0) & c1015(7) ;
		seg_scan <= not c1015;
	end if;

--if seg_a='1' then
--	segout<=x"ff";
--	segout_2<=x"ff";
--else
--end if;
	if c1015=x"04" then 	segout_2<="11000110";
	elsif c1015=x"40" then	segout	<="10110111";
	elsif c1015=x"80" then 	segout	<="11001111";
	else
		segout(7 downto 1)  <=seg_num(conv_integer(seg1));
		segout_2(7 downto 1)<=seg_num(conv_integer(seg2));
		segout(0)  <='0';
		segout_2(0)<='0';
	end if;
----------------------------------------------------------------------------
	--c1015
	--x"01" : 10000000	--x"02" : 01000000	--x"04" : 00100000	--x"08" : 00010000
	--x"10" : 00001000	--x"20" : 00000100	--x"40" : 00000010	--x"80" : 00000001
----------------------------------------------------------------------------
--	if c1015=x"02" then
--		segout_2(0)<='1';
--	else
--		segout_2(0)<='0';
--	end if;

end if;	
end if;

end process;
--========================================================================
BL  <= '1';
x<=CONV_INTEGER(add(6 DOWNTO 0));
y<=CONV_INTEGER(add(14 DOWNTO 7));
process(ck_LCD, nReset)          -- LCD
      variable delay_1         :integer range 0 to 25000000;                                                      	               	
      variable bit_cnt         :integer RANGE 0 TO 7 := 7;
      variable hi_lo           :integer range 0 to 1;
      variable address_start,address_end   : STD_LOGIC_VECTOR(14 DOWNTO 0); 	               	
      variable disp_color      : STD_LOGIC_VECTOR(5 DOWNTO 0); 	               	
      variable pos_x_start,pos_y_start :integer range 0 to 159;  
      variable pos_x,pos_y    :integer range 0 to 39;         
      variable pos_now              :integer range 0 to 20479;   	                  
      variable varl,cnt_number,cnt_number_max   :integer range 0 to 20;                                      
      variable cnt1           :integer range 0 to 99;                  
      variable bit_index   :integer range 0 to 16; 	               	
               
	begin	
      if(nReset ='0')then 
         RES <= '1';
         DC  <= '0';                              -- command
         CS  <= '1';
         SCL <= '1';                                     	                
         fsm <= 0;
         delay_1 :=0;
         address <= "0000000000000000";
                  
       else IF(ck_LCD'EVENT AND ck_LCD='1')then 
                      
     

--         if (event_S1 = '1') then                    -- �}�l�C��DEMO  
--                      
--            fsm <= 1;                        
--            DC  <= '0';                              -- �]���w�]��
--            CS  <= '1';
--            SCL <= '1';                                     	                
--            delay_1 :=0;
--            address <= "0000000000000000";
--            
--         elsif (event_S3 = '1') then                 -- �����C��DEMO
--            fsm <= 0;                        
--            DC  <= '0';                              -- �]���w�]��
--            CS  <= '1';
--            SCL <= '1';                                     	                
--            delay_1 :=0;
--            address <= "0000000000000000";
         
--         else
if (delay_1 )=0 then
            CASE fsm IS                                          
               when 0 =>   fsm <= 1;                           -- idle
                              
               when 1 =>                             -- �w��RESET, 0-2 
                        RES <= '1'; 
                        delay_1 :=25000;
                         fsm <= 2;                 
--                        if delay_1 >= 25000 then     -- 1ms = 40ns x 25000
--                           delay_1 :=0;                           
--                           fsm <= 2;
--                        else
--                           delay_1:=delay_1+1;                          
--                        end if;

               when 2 =>                             
                        RES <= '0';                  -- 1ms
                        delay_1 :=25000;
                        fsm <= 3;
--                        if delay_1 >= 25000 then                     
--                           delay_1 :=0;                           
--                           fsm <= 3;
--                        else
--                           delay_1:=delay_1+1;                          
--                        end if;

               when 3 =>                            
                        RES <= '1';                  -- 120ms
                        delay_1 :=3000000;
                        fsm <= 4;
--                        if delay_1 >= 3000000 then                
--                           delay_1 :=0;  
--                           fsm   <=  4;
--                           
--                        else
--                           delay_1:=delay_1+1;                          
--                        end if;               

               when 4 =>                                --start loop ,lcd��l�ƩR�O,�@85BYTES
                        if(address = "0000000001010101") then  
                           fsm        <= 5;                
                        else
                           fsm        <= 50;               
                           fsm_back   <=  4;            
                        end if;
                           
               when 5 =>   
                                    
                        delay_1 :=3000000;
                        fsm <= 6;                             -- ��l�ƫ᩵��    
--                        if delay_1 >= 3000000 then       -- 120ms                                         
--                           delay_1 :=0; 
--                           fsm     <= 6; 
--                        else
--                           delay_1:=delay_1+1;                          
--                        end if;

               when 6 =>                                -- idle   
--                        if (mode = 0) then
--                           fsm     <= 60; 
--                        elsif ((mode = 1) or (mode = 3)) then   
                           fsm     <= 10;   
--                        elsif (mode = 2) then   
--                           fsm     <= 110;                                                                                  
--                        end if;                                                                     
               
               when 10 =>                                ----------------------��s�e��,DISP_WINDOWS ,10-13     
                        address <= "0000000001001010";                     
                        fsm        <= 11;                

               when 11 =>                                --loop ,DISP_WINDOWS �R�O    
                        if(address = "0000000001010101") then  --�@11BYTES
                           add <= "000000000000000";
                           fsm        <= 12;                
                        else
                           fsm        <= 50;               
                           fsm_back   <= 11;            
                        end if;
                           
               when 12 =>                              -- start loop ,read ram                                 
                        hi_lo := 0;
                        we2  <= '0';
						if(add = 20480) then  fsm <= 10;LCD_t<=LCD_t+1;else add<=add+1;--fsm_back2;  -- ������s --                        a2   <= address(14 downto 0);               -- set address                                           
                        fsm  <= 13; end if;                       

               when 13 =>                              -- read ram                                 
                        if(hi_lo = 0)then              -- COLOR HI BYTE 
                                                       -- R - f800   G - 07e0  B - 001f 
                           RGB_data <= RGB(15 downto 8);
                                         
                              
                           
                              fsm        <= 40;               
                              fsm_back   <= 13;            
--                           end if;
                                                                                 
                        else                             --COLOR LO BYTE                         
                           RGB_data <=  RGB(7 downto 0);
                              
                           fsm        <= 40;  
                           fsm_back   <= 12;                                                     
                        end if;                      

--               when 20 =>                                    --write ram -�����M��,����,20-26
--                        address <= '0' & address_start;                     
--                        fsm     <= 21;
--
--               when 21 =>                                    
--                        a2   <= address(14 downto 0);        -- set address                                                                
--                        fsm  <= 22;
--                        
--               when 22 =>                                    -- set data
--                        di2  <= disp_color;                  
--                        fsm  <= 23; 
--                        
--               when 23 =>                                    -- write
--                        we2  <= '1';
--                        fsm  <= 24; 
--
--               when 24 =>                                    -- write
--                        we2  <= '0';
--                        fsm  <= 25; 
--
--               when 25 =>                                    -- address
--                        address <= address + "0000000000000001";                                                                
--                        fsm  <= 26; 
--                        
--               when 26 =>                                    -- address
--                        if(address = address_end) then       -- 128 * 160
--                           fsm        <= fsm_back;                
--                        else
--                           fsm        <= 21;               
--                        end if;                                    
                  

               when 40 =>                             --------------------------------- write data START,40-45 
                        DC  <= '1';    
                        fsm <= 41; 
               when 41 =>                             -- CS = 0              
                        CS  <= '0';
                        bit_cnt := 7;  
                        fsm <= 42;                       
               
               when 42 =>                             -- LOOP x 8 ,set data            
                        SDA <= RGB_data(bit_cnt); 
                        fsm <= 43;                      
                        
               when 43 =>                             -- CLK = 0 
                        SCL <= '0';                           
                        fsm <= 44;
                                              
               when 44 =>                             -- CLK = 1 
                        SCL <= '1';                           
                        bit_cnt := bit_cnt - 1;
                        
                        if bit_cnt >= 7 then
                           fsm <= 45;                      
                        else
                           fsm <= 42;                                           
                        end if;
                           
               when 45 =>                             -- CS = 1              
                        CS  <= '1';                     
                        if(hi_lo = 0)then
                           hi_lo := 1;
                        else
                           hi_lo := 0; 
                           address <= address + "0000000000000001";                          
                        end if;   
                        fsm <= fsm_back;                                                               

               when 50 =>                             -------------------------- write command START,50-55
                        DC  <= DC_data;    
                        fsm <= 51;                     
                        
               when 51 =>                             -- CS = 0              
                        CS  <= '0';
                        bit_cnt := 7;  
                        fsm <= 52;                       
               
               when 52 =>                             -- LOOP x 8 ,set data            
                        SDA <= data_out(bit_cnt); 
                        fsm <= 53;                      
                        
               when 53 =>                             -- CLK = 0 
                        SCL <= '0';                           
                        fsm <= 54;
                                              
               when 54 =>                             -- CLK = 1 
                        SCL <= '1';                           
                        bit_cnt := bit_cnt - 1;
                        
                        if bit_cnt >= 7 then
                           fsm <= 55;                      
                        else
                           fsm <= 52;                                           
                        end if;
                           
               when 55 =>                             -- CS = 1              
                        CS  <= '1';
                        address <= address + "0000000000000001"; 
                        fsm <= fsm_back;             

   ----------------------------------------------------------------------------       
               when 59 =>
                                       
                        delay_1 :=25000000;
                        fsm <=fsm_back2;                                 -- delay 1s
--                        if delay_1 >= 25000000 then                     
--                           delay_1 :=0;                           
--                           fsm <= fsm_back2;
--                        else
--                           delay_1:=delay_1+1;                          
--                        end if;
   ----------------------------------------------------------------------------  MODE = "00" ,�C��i��    
--               when 60 =>                                   -- 1 �ק�ϫ�    
--                        address_start := "000000000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "111111";          -- R - f800   G - 07e0  B - 001f                    
--                        fsm       <= 20;                   
--                        fsm_back  <= 61;                             
--
--               when 61 =>                                   --��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 62;   
--
--               when 62 =>                                   -- delay 1s  
--                        delay_1 :=0; 
--                        fsm       <= 59;                           
--                        fsm_back2 <= 63;
--                                
--               when 63 =>                                  -- 2 �ק�ϫ�                                                             
--                        address_start := "000000000000000";
--                        address_end   := "001100100000000";
--                        disp_color    := "000001";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 64;                             
--    
--               when 64 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 65;
--
--               when 65 =>                                  -- delay 1s  
--                        delay_1 :=0;    
--                        fsm       <= 59;                       
--                        fsm_back2 <= 66;
--
--               when 66 =>                                  -- 3 �ק�ϫ� 
--                        address_start := "000000000000000";
--                        address_end   := "001100100000000";
--                        disp_color    := "000010";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 67;
--
--               when 67 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 68;
--
--               when 68 =>                                  -- delay 1s  
--                        delay_1 :=0; 
--                        fsm       <= 59;                           
--                        fsm_back2 <= 69;
--               
--               when 69 =>                                  -- 4
--                        address_start := "000000000000000";
--                        address_end   := "001100100000000";
--                        disp_color    := "000011";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 70;
--
--               when 70 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 71;
--
--               when 71 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 72;           
--
--               when 72 =>                                  -- 5
--                        address_start := "001100100000000";
--                        address_end   := "011001000000000";
--                        disp_color    := "010000";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 73;
--
--               when 73 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 74;
--
--               when 74 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 75; 
--
--
--               when 75 =>                                  -- 6
--                        address_start := "001100100000000";
--                        address_end   := "011001000000000";
--                        disp_color    := "100000";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 76;
--
--               when 76 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 77;
--
--               when 77 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 78;
--
--               when 78 =>                                  -- 7
--                        address_start := "001100100000000";
--                        address_end   := "011001000000000";
--                        disp_color    := "110000";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 79;
--
--               when 79 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 80;
--
--               when 80 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 81;
--
--               when 81 =>                                  -- 8
--                        address_start := "011001000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "000100";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 82;
--
--               when 82 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 83;
--
--               when 83 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 84;
--
--               when 84 =>                                  -- 9
--                        address_start := "011001000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "001000";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 85;
--
--               when 85 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 86;
--
--               when 86 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 87;
--
--               when 87 =>                                  -- 10
--                        address_start := "011001000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "001100";         -- R"00"G"00"B"00"                   
--                        fsm       <= 20;                   
--                        fsm_back  <= 88;
--
--               when 88 =>                                  -- ��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 89;
--
--               when 89 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 90;
--
--               when 90 =>                                  -- delay 1s  
--                        delay_1 :=0;  
--                        fsm       <= 59;                          
--                        fsm_back2 <= 91;
--                        
--               when 91 =>                                  -- LOOP,���G
--                        address_start := "000000000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "111111";         -- R - f800   G - 07e0  B - 001f                    
--                        fsm       <= 20;                   
--                        fsm_back  <= 63;                              

   ----------------------------------------------------------------------------  MODE = "01" ,�զ���G
--               when 100 =>                                   -- 1 �ק�ϫ�    
--                        address_start := "000000000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "111100";          -- R - f800   G - 07e0  B - 001f                    
--                        fsm       <= 20;                   
--                        fsm_back  <= 101;                             
--
--               when 101 =>                                   --��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 102;   
--
--               when 102 =>                                   -- idle

   ----------------------------------------------------------------------------  MODE = "10" ,��ܤ�r �ϧ�, ���j�׼ƭ�
--               when 110 =>                                   -- �M���e��    
--                        address_start := "000000000000000";
--                        address_end   := "101000000000000";
--                        disp_color    := "111111";           -- ���G
--                        fsm       <= 20;                   
--                        fsm_back  <= 111;                             
--
--   ----------------------------------------------------------------------------�}�l�K�� 
--               when 111 =>                                   -- 1.��l���ܼ�   
--                        pos_x       := 0;
--                        pos_y       := 0;
--                        varl        := 0;                    -- ��ܤ�r�����
--                        cnt_number  := 0;                    -- �ثe��ܲĴX�Ӥ�r                        
--                        cnt_number_max := 9;                 -- �n��ܪ���r�ƶq   
--                        cnt1        := 0;                    -- 
--                        bit_index   := 15;                   -- 
--                        fsm         <= 113;   
--                                               
--               when 112 =>                                   -- 2.�]�w��ܤ�r & �K�Ϧ�m                    
--               	      if (cnt_number = 0) then             --   LOOP 112-119 
--                           varl := lx1;    
--                           if TSL2561_int > 20 then
--                              disp_color  := "000000";          -- ��r���C��,��                                                                                                       
--                              motor_dir <= '0';                  -- ���F����
--                           else
--                              disp_color  := "001100";          -- ��r���C��,��   
--                              motor_dir <= '1';                  -- ���F����
--                           end if;                              
--                           pos_x_start  := 20;
--                           pos_y_start  := 20;                
--                        elsif (cnt_number = 1)  then                            
--                           varl := lx2;    
--                           pos_x_start  := 36;
--                           pos_y_start  := 20;                                          
--                        elsif (cnt_number = 2)  then                            
--                           varl := lx3;
--                           pos_x_start  := 52;
--                           pos_y_start  := 20;                                          
--                        elsif (cnt_number = 3)  then                                                      
--                           varl := lx4;
--                           pos_x_start  := 68;                           
--                           pos_y_start  := 20; 
--                        elsif (cnt_number = 4)  then                                                      
--                           varl := lx5;
--                           pos_x_start  := 84;                           
--                           pos_y_start  := 20;                            
--                        elsif (cnt_number = 5)  then                                                      
--                           varl := 11;                       -- 'R'
--                           disp_color  := "000000";          -- ��r���C��,��
--                           pos_x_start  := 20;                           
--                           pos_y_start  := 60; 
--                        elsif (cnt_number = 6)  then                                                      
--                           varl := 12;                       -- 'T'
--                           disp_color  := "000000";          -- ��r���C��,��
--                           pos_x_start  := 36;                           
--                           pos_y_start  := 60;   
--                        elsif (cnt_number = 7)  then                                                      
--                           varl := 13;                       -- ':'
--                           disp_color  := "000000";          -- ��r���C��,��
--                           pos_x_start  := 52;                           
--                           pos_y_start  := 60;  
--                        elsif (cnt_number = 8)  then   
--                           if TSL2561_int > 20 then                                                   
--                              varl := 14;                       -- '���f��'
--                              disp_color  := "000000";          -- ��r���C��,��
--                           else
--                              varl := 15;                       -- '���f��'
--                              disp_color  := "110000";          -- ��r���C��,��                              
--                           end if;      
--                           pos_x_start  := 80;                           
--                           pos_y_start  := 60;                                                                                                                                                                                         
--                        end if;
--                        fsm       <= 113;                   
--                        
--               when 113 =>                                     -- 2.�]�wLCD��},�d��0 - (128*160-1)  ,111-115����8�I(1��BYTE)����Ƽg�J
--                        pos_now := pos_x_start + ((pos_y_start + pos_y) * 128) + pos_x;    
--                        pos_x   := pos_x + 1;
--                         
--                        fsm       <= 114;                   
--
--               when 114 =>                                     -- set address 
--                        a2   <= conv_std_logic_vector(pos_now,15);                                                                    
--                        fsm  <= 115;
--                        
--               when 115 =>                                     -- set data
--                        if(num_table(varl, cnt1)(bit_index) = '1') then                                                      
--                           di2  <= disp_color;                 --                              
--                        else
--                           di2  <= "111111";                                             
--                        end if;    
--                           
--                        fsm  <= 116; 
--                        
--               when 116 =>                                     -- write
--                        we2  <= '1';
--                        fsm  <= 117; 
--
--               when 117 =>                                     -- write
--                        we2  <= '0';
--                        
--                        if pos_x >= 16 then                    --�r��e��20
--                           pos_x := 0; 
--                           pos_y := pos_y + 1;                 --�r�鰪��40(40/8byte = 5)
--                        end if;
--                                                                           
--                        if(bit_index = 0) then
--                           bit_index := 15;
--                           fsm  <= 118; 
--                        else   
--                           bit_index   := bit_index - 1;                                             
--                           fsm  <= 113;                         
--                        end if;
--                                                
--               when 118 =>                                                               
--                           if cnt1 >= 15 then                  --�C�ӼƦr15��word(16bits)
--                              cnt1 := 0;
--                              fsm  <= 119; 
--                           else
--                              cnt1 := cnt1 + 1;                     
--                              fsm  <= 112; 
--                           end if;
--                        
--               when 119 =>                                    
--                        if (cnt_number < (cnt_number_max-1)) then  -- ��ܼƶq
--                           cnt_number := cnt_number + 1;           -- ����U�ӼƦr                                                                                 
--                           pos_x       := 0;
--                           pos_y       := 0;
--                           
--                           fsm       <= 113;      
--                        else
--                           cnt_number := 0;
--                           fsm       <= 120;                                
--                        end if;   
--               
--               when 120 =>                                   --��s�e��    
--                        fsm       <= 10;                   
--                        fsm_back2 <= 121;                  
--
--               when 121 =>                                  -- delay 1s , 1���s1�����  
--                        delay_1 :=0; 
--                        fsm       <= 59;                           
--                        fsm_back2 <= 110;
--               
               when others =>                          
                             
            END CASE;    
         
            
  

                  
                                        
	else delay_1 :=delay_1 -1;                             
    end if;
             end if; 
                      end if;  	   
	end process;
--=================================================================MOTOR_control--1
MOTOR_control1:process(nReset, ck_mot)           -- MOTOR-PWM
 	   variable scan_number    :integer range 0 to 9; 	 
   begin	
      if(nReset='0')then 	
         motor_out1 <= '0';
         motor_out2 <= '0';
         motor_pwm1 <= '0';
         scan_number := 0;
         
      elsif(ck_mot 'event and ck_mot ='1')then
         
--         if(mode_motor = 1) then                
 
             if(motor_dir1 = '0') then
               motor_out1 <= '1';                   --����
               motor_out2 <= '0';            
            else           
               motor_out1 <= '0';                   --����
               motor_out2 <= '1';                           
            end if;  
            
            if(scan_number >= 9) then 
               scan_number := 0;
            else      
               scan_number := scan_number + 1;                        
            end if;   
               
            if(motor_speed1 > scan_number) then 
               motor_pwm1 <= '1';
               --PWM1<='1';
            else      
               motor_pwm1 <= '0';
               --PWM1<='0';
            end if; 

--         elsif(mode_motor = 2) then                 --���t
--            motor_pwm1 <= '1';                   
            
          
                                                                
--         else
--            motor_out1 <= '0';
--            motor_out2 <= '0';
--            motor_pwm1 <= '0';
--            scan_number := 0;            
--               
--         end if;                         
                                    
      end if;   

   end process;
--=================================================================MOTOR_control--1
MOTOR_control2:process(nReset, ck_mot)           -- MOTOR-PWM
variable scan_number    :integer range 0 to 9; 	 
begin	
  if(nReset='0')then 	
	 motor_out3 <= '0';
	 motor_out4 <= '0';
	 motor_pwm2 <= '0';
	 scan_number := 0;
	 
  elsif(ck_mot 'event and ck_mot ='1')then
	 
--         if(mode_motor = 1) then                
 
		 if(motor_dir2 = '0') then
		   motor_out3 <= '1';                   --����
		   motor_out4 <= '0';            
		else           
		   motor_out3 <= '0';                   --����
		   motor_out4 <= '1';                           
		end if;  
		
		if(scan_number >= 9) then 
		   scan_number := 0;
		else      
		   scan_number := scan_number + 1;                        
		end if;   
		   
		if(motor_speed2 > scan_number) then 
		   motor_pwm2 <= '1';
		  -- PWM2<='1';
		else      
		   motor_pwm2 <= '0';
		 --  PWM2<='0';
		end if;                         
								
  end if;   

end process;
--===============================================================================RS232 to PC
topc:process(ck_1M) --press bt then sent dataT to pc
variable s:integer range 0 to 3;
variable t:integer range 0 to 51;
variable y:integer range 0 to 8;
variable x:integer range 0 to 7;--  0-1, 0-3, 0-7, 0-15, 0-31......
begin

if rising_edge(ck_1M) then
btt<=bt;
		if t = 0 then
		
			case s is
			
			when 0 =>
				if bt='1' and btt='0' then 
					
					s := 1;
					RSout <= '0'; 
					t := 25;
					y := 0;
				else 
					RSout <= '1';
				end if;
				
			when 1 =>
			
				if y = 8 then 
					y := 0;
					x := x+1;
					s := 2;
					RSout <= '1';
					t := 51;
				else 
					RSout <= dataT(x)(y); 
					t := 25;
					y := y+1;--tx datdR
				end if;
				
			when 2 =>
			
				if x = 0 then 
					s := 3;
				else 
					s := 1;
					RSout <= '0'; 
					t := 25;
				end if;
							 
			when 3 =>
			
				--if bt = '0'then 
					s := 0;t:=51;--t:=51;is the fast
				--end if;
				
			when others => null;
			end case;
		
	else t:=t-1;
	end if;
end if;
end process;
--====================================================================================
from_pc:process(ck_1M)	--recever pcdata to dataR

variable ib:std_logic;
variable y:integer range 0 to 8;
variable t:integer range 0 to 38 ;
variable x:integer range 0 to 1;--  0-1, 0-3, 0-7, 0-15, 0-31......
begin

if rising_edge(ck_1M) then

	if ib = '0' then 
		ib := not RSin;
		t := 38;
	else 
		if t = 0 then 
			if y = 8 then 
				y := 0;
				x := x+1;
				ib := '0';
				if x = 0 then 
					PcOkFlag <= not PcOkFlag;
				end if;--PcOkFlag is to main singal
			else 
				dataR(x)(y) <= RSin; 
				t := 25; 
				y := y+1;
			end if;
		 else 
			t := t-1;
		 end if;
	end if;
end if;
end process;
------------------------------------------------------------------------�s��w 
   u0:i2c_master        --SD178�X�� �Ҩϥ�IIC
   generic map 
   (
	  input_clk => 50_000_000,
	  bus_clk   => 10_000               --10_000
   )
   port map 
   (
	 clk       => ck,
	 reset_n   => sd178_nrst,
    
    ena       => sd178_ena, 
    addr      => "0100000",--sd178_addr
    
    rw        => sd178_rw, 
    data_wr   => sd178_data_wr,
    busy      => sd178_busy,
    data_rd   => sd178_data_rd, 
    ack_error => open,
    sda       => SD178_sda,
    scl       => SD178_scl
   );            

   u1:TSL2561
   port map(
         clk_50M => ck,
         nrst    => nReset,    
         
         sda       => TSL2561_sda,
         scl       => TSL2561_scl,
         
         TSL2561_data => TSL2561_data

           );

   u2:DHT11
   port map(
         clk_50M => ck,
         nrst    => nReset,    
         dat_bus => SHT11_PIN,
         HU      => HU_BUFF,
         TE      => TE_BUFF,                 
         error   => DHT11_error 

           );
 

   u9:cmd_rom           --��l�ƩR�O���
   port map 
   (
	 address   => address,
    data_out  => data_out,
    DC_data   => DC_data 
   );

--   u10:raminfr          --LCD ��ܸ�ƼȦsRAM
--   generic map 
--	 (
--		  bits        => 6,
--		  addr_bits   => 15              
--	 )            
--   port map(      
--               clk     => ck,       
--	            we      => we2,
--               a       => a2,
--               di      => di2,
--               do      => do2   
--            );
--          
                 
end beh;